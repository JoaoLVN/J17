// [[Joe - joao.euu@gmail.com]]

module J17 ();

endmodule //
