// [[Joe - joao.euu@gmail.com]]

module J17 ( input clk ,output [31:0] result,output [31:0]instruct, output [31:0]progcount,output [3:0]alucd, output [2:0] o1,output [20:0] o2,output im);

 wire [31:0]PC;
 wire[31:0]instruction;

 wire [3:0] alucode;
 wire [2:0] op1;
 wire [20:0] op2;
 wire [3:0] pcControl;
 wire flag;
 wire flag1;
 wire imControl;
 wire writecode;
 wire [1:0] stackSelect;

 assign instruct=instruction;
 assign progcount=PC;
 assign alucd=alucode;
 assign o1=op1;
 assign o2=op2;
 assign im=imControl;


 IF InstructionFetch(
 .clock(clk),
 .pc(PC),
 .out(instruction)
 );

 UC ControlUnit(
 .clock(clk),
 .instruction(instruction),
 .alucode(alucode),
 .op1(op1),
 .op2(op2),
 .imControl(imControl),
 .writecode(writecode),
 .pcControl(pcControl),
 .flag(flag),
 .flag1(flag1),
 .stackSelect(stackSelect),
	);
DP DataPath(
  .clock(clk),
  .alucode(alucode),
  .flag(flag),
  .flag1(flag1),
  .op1(op1),
  .op2(op2),
  .imControl(imControl),
  .pcControl(pcControl),
  .writecode(writecode),
  .stackSelect(stackSelect),
  .PC(PC),
  .result(result)
  );



endmodule //
