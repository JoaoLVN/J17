// [[Joe - joao.euu@gmail.com]]

module ControlUnit ();

endmodule 
